Name: Sanduri Ashok Kumar
ID: CT12DS2126
Domain:vlsi
Duration: AUGUST 5th to OCTOBER 5th 2024

Overview of the Project

Project: Digital Design Verification

Heading: Finite State Machine (FSM) Design and Testbench

Key Activities:

- Designed and implemented a Finite State Machine (FSM) module in Verilog
- Created a testbench to verify the functionality of the FSM module
- Simulated the testbench using Xilinx Vivado Simulator

Technology:

- Digital Design
- Verilog HDL
- Finite State Machines

Tools Used:

- Xilinx Vivado Simulator
- Verilog Compiler

